kah704@quser31.quest.it.northwestern.edu.183989:1680277453